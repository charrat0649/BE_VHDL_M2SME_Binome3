  --Example instantiation for system 'RAMZI'
  RAMZI_inst : RAMZI
    port map(
      clk_adc_from_the_verin_test_0 => clk_adc_from_the_verin_test_0,
      cs_n_from_the_verin_test_0 => cs_n_from_the_verin_test_0,
      done_probe_from_the_avalon_txd_0 => done_probe_from_the_avalon_txd_0,
      internal_reset_from_the_gestion_anemometre_0 => internal_reset_from_the_gestion_anemometre_0,
      ledBabord_from_the_avalon_gestion_bp_0 => ledBabord_from_the_avalon_gestion_bp_0,
      ledSTBY_from_the_avalon_gestion_bp_0 => ledSTBY_from_the_avalon_gestion_bp_0,
      ledTribord_from_the_avalon_gestion_bp_0 => ledTribord_from_the_avalon_gestion_bp_0,
      out_bip_from_the_avalon_gestion_bp_0 => out_bip_from_the_avalon_gestion_bp_0,
      out_port_from_the_sortie => out_port_from_the_sortie,
      out_pwm_from_the_avalon_pwm_0 => out_pwm_from_the_avalon_pwm_0,
      out_pwm_from_the_verin_test_0 => out_pwm_from_the_verin_test_0,
      out_sens_from_the_verin_test_0 => out_sens_from_the_verin_test_0,
      readdata_from_the_avalon_txd_0 => readdata_from_the_avalon_txd_0,
      txd_from_the_avalon_txd_0 => txd_from_the_avalon_txd_0,
      BP_Babord_to_the_avalon_gestion_bp_0 => BP_Babord_to_the_avalon_gestion_bp_0,
      BP_STBY_to_the_avalon_gestion_bp_0 => BP_STBY_to_the_avalon_gestion_bp_0,
      BP_Tribord_to_the_avalon_gestion_bp_0 => BP_Tribord_to_the_avalon_gestion_bp_0,
      clk_0 => clk_0,
      data_in_to_the_verin_test_0 => data_in_to_the_verin_test_0,
      in_freq_anemometre_to_the_gestion_anemometre_0 => in_freq_anemometre_to_the_gestion_anemometre_0,
      in_port_to_the_entree => in_port_to_the_entree,
      in_pwm_compas_to_the_avalon_compas_0 => in_pwm_compas_to_the_avalon_compas_0,
      reset_n => reset_n
    );


